
module Fonts(FontSelect,PosFila,Fila);

input [4:0] FontSelect;
input [3:0] PosFila;
output [15:0] Fila;

reg[15:0] Fila;

always@(FontSelect or PosFila) 
	case ({FontSelect,PosFila})
	//CERO
		9'b000000000:  Fila = 16'b0000000000000000;
		9'b000000001:  Fila = 16'b0000000000000000;
		9'b000000010:  Fila = 16'b0000011111100000;
		9'b000000011:  Fila = 16'b0000110000110000;
		9'b000000100:  Fila = 16'b0001100000011000;
		9'b000000101:  Fila = 16'b0001100000011000;
		9'b000000110:  Fila = 16'b0001100000011000;
		9'b000000111:  Fila = 16'b0001100000011000;
		9'b000001000:  Fila = 16'b0001100000011000;
		9'b000001001:  Fila = 16'b0001100000011000;
		9'b000001010:  Fila = 16'b0001100000011000;
		9'b000001011:  Fila = 16'b0001100000011000;
		9'b000001100:  Fila = 16'b0000110000110000;
		9'b000001101:  Fila = 16'b0000011111100000;
		9'b000001110:  Fila = 16'b0000000000000000;
		9'b000001111:  Fila = 16'b0000000000000000;
	//UNO
		9'b000010000: Fila =  16'b0000000000000000;
		9'b000010001: Fila =  16'b0000000000000000;
		9'b000010010: Fila =  16'b0000000000000000;
		9'b000010011: Fila =  16'b0000000110000000;
		9'b000010100: Fila =  16'b0000001110000000;
		9'b000010101: Fila =  16'b0000111110000000;
		9'b000010110: Fila =  16'b0000000110000000;
		9'b000010111: Fila =  16'b0000000110000000;
		9'b000011000: Fila =  16'b0000000110000000;
		9'b000011001: Fila =  16'b0000000110000000;
		9'b000011010: Fila =  16'b0000000110000000;
		9'b000011011: Fila =  16'b0000000110000000;
		9'b000011100: Fila =  16'b0000000110000000;
		9'b000011101: Fila =  16'b0000111111110000;
		9'b000011110: Fila =  16'b0000000000000000;
		9'b000011111: Fila =  16'b0000000000000000;
	//DOS
		9'b000100000: Fila =  16'b0000000000000000;
		9'b000100001: Fila =  16'b0000000000000000;
		9'b000100010: Fila =  16'b0000011111000000;
		9'b000100011: Fila =  16'b0000110001100000;
		9'b000100100: Fila =  16'b0001100000110000;
		9'b000100101: Fila =  16'b0001100000110000;
		9'b000100110: Fila =  16'b0000000001100000;
		9'b000100111: Fila =  16'b0000000011000000;
		9'b000101000: Fila =  16'b0000000110000000;
		9'b000101001: Fila =  16'b0000001100000000;
		9'b000101010: Fila =  16'b0000011000000000;
		9'b000101011: Fila =  16'b0000110000000000;
		9'b000101100: Fila =  16'b0001100000000000;
		9'b000101101: Fila =  16'b0001111111110000;
		9'b000101110: Fila =  16'b0000000000000000;
		9'b000101111: Fila =  16'b0000000000000000;
	//TRES
		9'b000110000: Fila =  16'b0000000000000000;
		9'b000110001: Fila =  16'b0000000000000000;
		9'b000110010: Fila =  16'b0000011111100000;
		9'b000110011: Fila =  16'b0000110000110000;
		9'b000110100: Fila =  16'b0001100000011000;
		9'b000110101: Fila =  16'b0000000000011000;
		9'b000110110: Fila =  16'b0000000000110000;
		9'b000110111: Fila =  16'b0000001111110000;
		9'b000111000: Fila =  16'b0000001111110000;
		9'b000111001: Fila =  16'b0000000000110000;
		9'b000111010: Fila =  16'b0000000000011000;
		9'b000111011: Fila =  16'b0001100000011000;
		9'b000111100: Fila =  16'b0000110000110000;
		9'b000111101: Fila =  16'b0000011111100000;
		9'b000111110: Fila =  16'b0000000000000000;
		9'b000111111: Fila =  16'b0000000000000000;
	//CUATRO
		9'b001000000: Fila =  16'b0000000000000000;
		9'b001000001: Fila =  16'b0000000000000000;
		9'b001000010: Fila =  16'b0001100001100000;
		9'b001000011: Fila =  16'b0001100001100000;
		9'b001000100: Fila =  16'b0001100001100000;
		9'b001000101: Fila =  16'b0001100001100000;
		9'b001000110: Fila =  16'b0001100001100000;
		9'b001000111: Fila =  16'b0001100001100000;
		9'b001001000: Fila =  16'b0001111111111000;
		9'b001001001: Fila =  16'b0000000001100000;
		9'b001001010: Fila =  16'b0000000001100000;
		9'b001001011: Fila =  16'b0000000001100000;
		9'b001001100: Fila =  16'b0000000001100000;
		9'b001001101: Fila =  16'b0000000001100000;
		9'b001001110: Fila =  16'b0000000000000000;
		9'b001001111: Fila =  16'b0000000000000000;
	//CINCO
		9'b001010000: Fila =  16'b0000000000000000;
		9'b001010001: Fila =  16'b0000000000000000;
		9'b001010010: Fila =  16'b0001111111111000;
		9'b001010011: Fila =  16'b0001100000000000;
		9'b001010100: Fila =  16'b0001100000000000;
		9'b001010101: Fila =  16'b0001100000000000;
		9'b001010110: Fila =  16'b0001100000000000;
		9'b001010111: Fila =  16'b0001111111100000;
		9'b001011000: Fila =  16'b0000000000110000;
		9'b001011001: Fila =  16'b0000000000011000;
		9'b001011010: Fila =  16'b0000000000011000;
		9'b001011011: Fila =  16'b0000000000011000;
		9'b001011100: Fila =  16'b0000000000110000;
		9'b001011101: Fila =  16'b0001111111100000;
		9'b001011110: Fila =  16'b0000000000000000;
		9'b001011111: Fila =  16'b0000000000000000;
	//SEIS
		9'b001100000: Fila =  16'b0000000000000000;
		9'b001100001: Fila =  16'b0000000000000000;
		9'b001100010: Fila =  16'b0000111111110000;
		9'b001100011: Fila =  16'b0001100000011000;
		9'b001100100: Fila =  16'b0001100000000000;
		9'b001100101: Fila =  16'b0001100000000000;
		9'b001100110: Fila =  16'b0001100000000000;
		9'b001100111: Fila =  16'b0001100000000000;
		9'b001101000: Fila =  16'b0001111111110000;
		9'b001101001: Fila =  16'b0001100000011000;
		9'b001101010: Fila =  16'b0001100000011000;
		9'b001101011: Fila =  16'b0001100000011000;
		9'b001101100: Fila =  16'b0001100000011000;
		9'b001101101: Fila =  16'b0000111111110000;
		9'b001101110: Fila =  16'b0000000000000000;
		9'b001101111: Fila =  16'b0000000000000000;
	//SIETE
		9'b001110000: Fila =  16'b0000000000000000;
		9'b001110001: Fila =  16'b0000000000000000;
		9'b001110010: Fila =  16'b0001111111111000;
		9'b001110011: Fila =  16'b0000000000011000;
		9'b001110100: Fila =  16'b0000000000011000;
		9'b001110101: Fila =  16'b0000000000011000;
		9'b001110110: Fila =  16'b0000000000110000;
		9'b001110111: Fila =  16'b0000000001100000;
		9'b001111000: Fila =  16'b0000000011000000;
		9'b001111001: Fila =  16'b0000000110000000;
		9'b001111010: Fila =  16'b0000000110000000;
		9'b001111011: Fila =  16'b0000000110000000;
		9'b001111100: Fila =  16'b0000000110000000;
		9'b001111101: Fila =  16'b0000000110000000;
		9'b001111110: Fila =  16'b0000000000000000;
		9'b001111111: Fila =  16'b0000000000000000;
	//OCHO
		9'b010000000: Fila =  16'b0000000000000000;
		9'b010000001: Fila =  16'b0000000000000000;
		9'b010000010: Fila =  16'b0000011111100000;
		9'b010000011: Fila =  16'b0000110000110000;
		9'b010000100: Fila =  16'b0001100000011000;
		9'b010000101: Fila =  16'b0001100000011000;
		9'b010000110: Fila =  16'b0000110000110000;
		9'b010000111: Fila =  16'b0000011111100000;
		9'b010001000: Fila =  16'b0000011111100000;
		9'b010001001: Fila =  16'b0000110000110000;
		9'b010001010: Fila =  16'b0001100000011000;
		9'b010001011: Fila =  16'b0001100000011000;
		9'b010001100: Fila =  16'b0000110000110000;
		9'b010001101: Fila =  16'b0000011111100000;
		9'b010001110: Fila =  16'b0000000000000000;
		9'b010001111: Fila =  16'b0000000000000000;
	//NUEVE
		9'b010010000: Fila =  16'b0000000000000000;
		9'b010010001: Fila =  16'b0000000000000000;
		9'b010010010: Fila =  16'b0000011111100000;
		9'b010010011: Fila =  16'b0000110000110000;
		9'b010010100: Fila =  16'b0001100000011000;
		9'b010010101: Fila =  16'b0001100000011000;
		9'b010010110: Fila =  16'b0001100000011000;
		9'b010010111: Fila =  16'b0000110000011000;
		9'b010011000: Fila =  16'b0000011111111000;
		9'b010011001: Fila =  16'b0000000000011000;
		9'b010011010: Fila =  16'b0000000000011000;
		9'b010011011: Fila =  16'b0000000000011000;
		9'b010011100: Fila =  16'b0000000000110000;
		9'b010011101: Fila =  16'b0000111111100000;
		9'b010011110: Fila =  16'b0000000000000000;
		9'b010011111: Fila =  16'b0000000000000000;
	//A
		9'b010100000: Fila =  16'b0000000000000000;
		9'b010100001: Fila =  16'b0000000000000000;
		9'b010100010: Fila =  16'b0000011111100000;
		9'b010100011: Fila =  16'b0000110000110000;
		9'b010100100: Fila =  16'b0001100000011000;
		9'b010100101: Fila =  16'b0001100000011000;
		9'b010100110: Fila =  16'b0001100000011000;
		9'b010100111: Fila =  16'b0001100000011000;
		9'b010101000: Fila =  16'b0001111111111000;
		9'b010101001: Fila =  16'b0001100000011000;
		9'b010101010: Fila =  16'b0001100000011000;
		9'b010101011: Fila =  16'b0001100000011000;
		9'b010101100: Fila =  16'b0001100000011000;
		9'b010101101: Fila =  16'b0001100000011000;
		9'b010101110: Fila =  16'b0000000000000000;
		9'b010101111: Fila =  16'b0000000000000000;
	//B
		9'b010110000: Fila =  16'b0000000000000000;
		9'b010110001: Fila =  16'b0000000000000000;
		9'b010110010: Fila =  16'b0001111111100000;
		9'b010110011: Fila =  16'b0001100000110000;
		9'b010110100: Fila =  16'b0001100000011000;
		9'b010110101: Fila =  16'b0001100000011000;
		9'b010110110: Fila =  16'b0001100000110000;
		9'b010110111: Fila =  16'b0001111111100000;
		9'b010111000: Fila =  16'b0001111111100000;
		9'b010111001: Fila =  16'b0001100000110000;
		9'b010111010: Fila =  16'b0001100000011000;
		9'b010111011: Fila =  16'b0001100000011000;
		9'b010111100: Fila =  16'b0001100000110000;
		9'b010111101: Fila =  16'b0001111111100000;
		9'b010111110: Fila =  16'b0000000000000000;
		9'b010111111: Fila =  16'b0000000000000000;
	//C
		9'b011000000: Fila =  16'b0000000000000000;
		9'b011000001: Fila =  16'b0000000000000000;
		9'b011000010: Fila =  16'b0000111111110000;
		9'b011000011: Fila =  16'b0001100000011000;
		9'b011000100: Fila =  16'b0001100000011000;
		9'b011000101: Fila =  16'b0001100000000000;
		9'b011000110: Fila =  16'b0001100000000000;
		9'b011000111: Fila =  16'b0001100000000000;
		9'b011001000: Fila =  16'b0001100000000000;
		9'b011001001: Fila =  16'b0001100000000000;
		9'b011001010: Fila =  16'b0001100000000000;
		9'b011001011: Fila =  16'b0001100000011000;
		9'b011001100: Fila =  16'b0001100000011000;
		9'b011001101: Fila =  16'b0000111111110000;
		9'b011001110: Fila =  16'b0000000000000000;
		9'b011001111: Fila =  16'b0000000000000000;
	//D
		9'b011010000: Fila =  16'b0000000000000000;
		9'b011010001: Fila =  16'b0000000000000000;
		9'b011010010: Fila =  16'b0001111111100000;
		9'b011010011: Fila =  16'b0001100000110000;
		9'b011010100: Fila =  16'b0001100000011000;
		9'b011010101: Fila =  16'b0001100000011000;
		9'b011010110: Fila =  16'b0001100000011000;
		9'b011010111: Fila =  16'b0001100000011000;
		9'b011011000: Fila =  16'b0001100000011000;
		9'b011011001: Fila =  16'b0001100000011000;
		9'b011011010: Fila =  16'b0001100000011000;
		9'b011011011: Fila =  16'b0001100000011000;
		9'b011011100: Fila =  16'b0001100000110000;
		9'b011011101: Fila =  16'b0001111111100000;
		9'b011011110: Fila =  16'b0000000000000000;
		9'b011011111: Fila =  16'b0000000000000000;
	//E
		9'b011100000: Fila =  16'b0000000000000000;
		9'b011100001: Fila =  16'b0000000000000000;
		9'b011100010: Fila =  16'b0001111111111000;
		9'b011100011: Fila =  16'b0001100000000000;
		9'b011100100: Fila =  16'b0001100000000000;
		9'b011100101: Fila =  16'b0001100000000000;
		9'b011100110: Fila =  16'b0001100000000000;
		9'b011100111: Fila =  16'b0001100000000000;
		9'b011101000: Fila =  16'b0001111111100000;
		9'b011101001: Fila =  16'b0001100000000000;
		9'b011101010: Fila =  16'b0001100000000000;
		9'b011101011: Fila =  16'b0001100000000000;
		9'b011101100: Fila =  16'b0001100000000000;
		9'b011101101: Fila =  16'b0001111111111000;
		9'b011101110: Fila =  16'b0000000000000000;
		9'b011101111: Fila =  16'b0000000000000000;
	//F
		9'b011110000: Fila =  16'b0000000000000000;
		9'b011110001: Fila =  16'b0000000000000000;
		9'b011110010: Fila =  16'b0001111111111000;
		9'b011110011: Fila =  16'b0001100000000000;
		9'b011110100: Fila =  16'b0001100000000000;
		9'b011110101: Fila =  16'b0001100000000000;
		9'b011110110: Fila =  16'b0001100000000000;
		9'b011110111: Fila =  16'b0001100000000000;
		9'b011111000: Fila =  16'b0001111111000000;
		9'b011111001: Fila =  16'b0001100000000000;
		9'b011111010: Fila =  16'b0001100000000000;
		9'b011111011: Fila =  16'b0001100000000000;
		9'b011111100: Fila =  16'b0001100000000000;
		9'b011111101: Fila =  16'b0001100000000000;
		9'b011111110: Fila =  16'b0000000000000000;
		9'b011111111: Fila =  16'b0000000000000000;
	//SUMA
		9'b100000000: Fila =  16'b0000000000000000;
		9'b100000001: Fila =  16'b0000000110000000;
		9'b100000010: Fila =  16'b0000000110000000;
		9'b100000011: Fila =  16'b0000000110000000;
		9'b100000100: Fila =  16'b0000000110000000;
		9'b100000101: Fila =  16'b0000000110000000;
		9'b100000110: Fila =  16'b0000000110000000;
		9'b100000111: Fila =  16'b0111111111111110;
		9'b100001000: Fila =  16'b0111111111111110;
		9'b100001001: Fila =  16'b0000000110000000;
		9'b100001010: Fila =  16'b0000000110000000;
		9'b100001011: Fila =  16'b0000000110000000;
		9'b100001100: Fila =  16'b0000000110000000;
		9'b100001101: Fila =  16'b0000000110000000;
		9'b100001110: Fila =  16'b0000000110000000;
		9'b100001111: Fila =  16'b0000000000000000;
	//RESTA
		9'b100010000: Fila =  16'b0000000000000000;
		9'b100010001: Fila =  16'b0000000000000000;
		9'b100010010: Fila =  16'b0000000000000000;
		9'b100010011: Fila =  16'b0000000000000000;
		9'b100010100: Fila =  16'b0000000000000000;
		9'b100010101: Fila =  16'b0000000000000000;
		9'b100010110: Fila =  16'b0000000000000000;
		9'b100010111: Fila =  16'b0111111111111110;
		9'b100011000: Fila =  16'b0111111111111110;
		9'b100011001: Fila =  16'b0000000000000000;
		9'b100011010: Fila =  16'b0000000000000000;
		9'b100011011: Fila =  16'b0000000000000000;
		9'b100011100: Fila =  16'b0000000000000000;
		9'b100011101: Fila =  16'b0000000000000000;
		9'b100011110: Fila =  16'b0000000000000000;
		9'b100011111: Fila =  16'b0000000000000000;
	//MULTIPLICACION
		9'b100100000: Fila =  16'b0000000000000000;
		9'b100100001: Fila =  16'b0000000000000000;
		9'b100100010: Fila =  16'b0110000000000110;
		9'b100100011: Fila =  16'b0011000000001100;
		9'b100100100: Fila =  16'b0001100000011000;
		9'b100100101: Fila =  16'b0000110000110000;
		9'b100100110: Fila =  16'b0000011001100000;
		9'b100100111: Fila =  16'b0000001111000000;
		9'b100101000: Fila =  16'b0000001111000000;
		9'b100101001: Fila =  16'b0000011001100000;
		9'b100101010: Fila =  16'b0000110000110000;
		9'b100101011: Fila =  16'b0001100000011000;
		9'b100101100: Fila =  16'b0011000000001100;
		9'b100101101: Fila =  16'b0110000000000110;
		9'b100101110: Fila =  16'b0000000000000000;
		9'b100101111: Fila =  16'b0000000000000000;
	//DIVISION//19
		9'b100110000: Fila = 16'b0000000000000000;
		9'b100110001: Fila = 16'b0000000000000000;
		9'b100110010: Fila = 16'b0000000000000000;
		9'b100110011: Fila = 16'b0000000000000000;
		9'b100110100: Fila = 16'b0000000001110000;
		9'b100110101: Fila = 16'b0000000011100000;
		9'b100110110: Fila = 16'b0000000111000000;
		9'b100110111: Fila = 16'b0000001110000000;
		9'b100111000: Fila = 16'b0000011100000000;
		9'b100111001: Fila = 16'b0000111000000000;
		9'b100111010: Fila = 16'b0001110000000000;
		9'b100111011: Fila = 16'b0011100000000000;
		9'b100111100: Fila = 16'b0111000000000000;
		9'b100111101: Fila = 16'b0000000000000000;
		9'b100111110: Fila = 16'b0000000000000000;
		9'b100111111: Fila = 16'b0000000000000000;
	//RAIZ /20
		9'b101000000: Fila =  16'b0000000000000000;
		9'b101000001: Fila =  16'b0001111111111110;
		9'b101000010: Fila =  16'b0001111111111110;
		9'b101000011: Fila =  16'b0001100000000000;
		9'b101000100: Fila =  16'b0001100000000000;
		9'b101000101: Fila =  16'b0001100000000000;
		9'b101000110: Fila =  16'b0001100000000000;
		9'b101000111: Fila =  16'b0001100000000000;
		9'b101001000: Fila =  16'b0001100000000000;
		9'b101001001: Fila =  16'b0001100000000000;
		9'b101001010: Fila =  16'b1111100000000000;
		9'b101001011: Fila =  16'b0111100000000000;
		9'b101001100: Fila =  16'b0111100000000000;
		9'b101001101: Fila =  16'b0011100000000000;
		9'b101001110: Fila =  16'b0001100000000000;
		9'b101001111: Fila =  16'b0000000000000000;
	//BORRAR /21
		9'b101010000: Fila =  16'b0000000000000000;
		9'b101010001: Fila =  16'b0000000000000000;
		9'b101010010: Fila =  16'b0000000000000000;
		9'b101010011: Fila =  16'b0000010000000000;
		9'b101010100: Fila =  16'b0000110000000000;
		9'b101010101: Fila =  16'b0001110000000000;
		9'b101010110: Fila =  16'b0011110000000000;
		9'b101010111: Fila =  16'b0111111111111110;
		9'b101011000: Fila =  16'b0111111111111110;
		9'b101011001: Fila =  16'b0011110000000000;
		9'b101011010: Fila =  16'b0001110000000000;
		9'b101011011: Fila =  16'b0000110000000000;
		9'b101011100: Fila =  16'b0000010000000000;
		9'b101011101: Fila =  16'b0000000000000000;
		9'b101011110: Fila =  16'b0000000000000000;
		9'b101011111: Fila =  16'b0000000000000000;
	//IGUAL /22
		9'b101100000: Fila =  16'b0000000000000000;
		9'b101100001: Fila =  16'b0000000000000000;
		9'b101100010: Fila =  16'b0111111111111110;
		9'b101100011: Fila =  16'b0111111111111110;
		9'b101100100: Fila =  16'b0000000000000000;
		9'b101100101: Fila =  16'b0000000000000000;
		9'b101100110: Fila =  16'b0000000000000000;
		9'b101100111: Fila =  16'b0000000000000000;
		9'b101101000: Fila =  16'b0000000000000000;
		9'b101101001: Fila =  16'b0000000000000000;
		9'b101101010: Fila =  16'b0000000000000000;
		9'b101101011: Fila =  16'b0000000000000000;
		9'b101101100: Fila =  16'b0111111111111110;
		9'b101101101: Fila =  16'b0111111111111110;
		9'b101101110: Fila =  16'b0000000000000000;
		9'b101101111: Fila =  16'b0000000000000000;	
	//AC /23
		9'b101110000: Fila =  16'b0000000000000000;
		9'b101110001: Fila =  16'b0001100001111110;
		9'b101110010: Fila =  16'b0010010001000000;
		9'b101110011: Fila =  16'b0100001001000000;
		9'b101110100: Fila =  16'b0100001001000000;
		9'b101110101: Fila =  16'b0100001001000000;
		9'b101110110: Fila =  16'b0100001001000000;
		9'b101110111: Fila =  16'b0100001001000000;
		9'b101111000: Fila =  16'b0111111001000000;
		9'b101111001: Fila =  16'b0100001001000000;
		9'b101111010: Fila =  16'b0100001001000000;
		9'b101111011: Fila =  16'b0100001001000000;
		9'b101111100: Fila =  16'b0100001001000000;
		9'b101111101: Fila =  16'b0100001001000000;
		9'b101111110: Fila =  16'b0100001001111110;
		9'b101111111: Fila =  16'b0000000000000000;
		
	//VACIO /24
		9'b110000000: Fila =  16'b0000000000000000;
		9'b110000001: Fila =  16'b0000000000000000;
		9'b110000010: Fila =  16'b0000000000000000;
		9'b110000011: Fila =  16'b0000000000000000;
		9'b110000100: Fila =  16'b0000000000000000;
		9'b110000101: Fila =  16'b0000000000000000;
		9'b110000110: Fila =  16'b0000000000000000;
		9'b110000111: Fila =  16'b0000000000000000;
		9'b110001000: Fila =  16'b0000000000000000;
		9'b110000000: Fila =  16'b0000000000000000;
		9'b110001001: Fila =  16'b0000000000000000;
		9'b110001010: Fila =  16'b0000000000000000;
		9'b110001011: Fila =  16'b0000000000000000;
		9'b110001100: Fila =  16'b0000000000000000;
		9'b110001101: Fila =  16'b0000000000000000;
		9'b110001110: Fila =  16'b0000000000000000;
		9'b110001111: Fila =  16'b0000000000000000;
	//PUNTO  /25
		9'b110010000: Fila = 16'b0000000000000000;
		9'b110010001: Fila = 16'b0000000000000000;
		9'b110010010: Fila = 16'b0000000000000000;
		9'b110010011: Fila = 16'b0000000000000000;
		9'b110010100: Fila = 16'b0000000000000000;
		9'b110010101: Fila = 16'b0000000000000000;
		9'b110010110: Fila = 16'b0000000000000000;
		9'b110010111: Fila = 16'b0000000000000000;
		9'b110011000: Fila = 16'b0000000000000000;
		9'b110011001: Fila = 16'b0000011111000000;
		9'b110011010: Fila = 16'b0000111111100000;
		9'b110011011: Fila = 16'b0000111111100000;
		9'b110011100: Fila = 16'b0000111111100000;
		9'b110011101: Fila = 16'b0000011111000000;
		9'b110011110: Fila = 16'b0000000000000000;
		9'b110011111: Fila = 16'b0000000000000000;
		
		default Fila =  16'b0000000000000000;
	endcase
endmodule
					