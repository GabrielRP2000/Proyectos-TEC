
module DegoBorde(X,Y,POS,Borde);

input [4:0] X;
input [3:0] Y;
input [4:0] POS;
output reg Borde;
//????? ?????????????????????
always@(X or Y or POS)
	casez({X,Y,POS})
		14'b00000?????????: Borde = 1'b1; //BORDE IZQUIERDA
		14'b?????0000?????: Borde = 1'b1; //BORDE ARRIBA
		14'b01001?????????: Borde = 1'b1; //BORDE DERECHA
		14'b?????0101?????: Borde = 1'b1; //BORDE ABAJO
		
		14'b?????0010?????: Borde = 1'b1; //1ER FILA
		14'b?????0011?????: Borde = 1'b1; //2DA FILA
		14'b?????0100?????: Borde = 1'b1;	//3RA FILA
//		13'b?????0101?????: Borde = 1'b1;	//4TA FILA
//		13'b?????0110?????: Borde = 1'b1; //5TA FILA

		14'b11111?????????: Borde = 1'b0;	//PRED X
//		13'b?????1000?????: Borde = 1'b0;	//PRED Y

		14'b000010001?????: Borde = 1'b0; 
		14'b000011111?????: Borde = 1'b1;   //1ER COLUMNA
//		3'b000011111??????????????????????????: Borde = 1'b1;
//		3'b000011111?????: Borde = 1'b1;
		
		14'b000100001?????: Borde = 1'b0; 
		14'b000101111?????: Borde = 1'b1;  
//		3'b000101111??????????????????????????: Borde = 1'b1;	//2DA COLUMNA
//		3'b000101111??????????????????????????: Borde = 1'b1;
		
		14'b000110001?????: Borde = 1'b0; 
		14'b000111111?????: Borde = 1'b1;  //3ER COLUMNA
//		3'b000111111?????: Borde = 1'b1;
//		3'b000111111?????: Borde = 1'b1;
		
		14'b001000001?????: Borde = 1'b0; 
		14'b001001111?????: Borde = 1'b1;  
//		3'b001001111?????: Borde = 1'b1;	//4TA COLUMNA
//		3'b001001111?????: Borde = 1'b1;
		
		14'b001010001?????: Borde = 1'b0; 
		14'b001011111?????: Borde = 1'b1;   //5TA COLUMNA
//		3'b001011111?????: Borde = 1'b1;
//		3'b001011111?????: Borde = 1'b1;
		
		14'b001100001?????: Borde = 1'b0; 
		14'b001101111?????: Borde = 1'b1;  
//		3'b001101111?????: Borde = 1'b1;	//6MA COLUMNA
//		3'b001101111?????: Borde = 1'b1;

		14'b001110001?????: Borde = 1'b0; 
		14'b001111111?????: Borde = 1'b1;  //7VA COLUMNA
//		3'b001111111?????: Borde = 1'b1;
//		3'b001111111?????: Borde = 1'b1;

		14'b010000001?????: Borde = 1'b0; 
		14'b010001111?????: Borde = 1'b1;  
//		3'b010001111?????: Borde = 1'b1;	//8VA COLUMNA
//		3'b010001111?????: Borde = 1'b1;
		
		
		14'b01010011010100: Borde = 1'b1; //0
		14'b01011011010101: Borde = 1'b1; //1
		14'b01100011010110: Borde = 1'b1; //2
		14'b01101011010111: Borde = 1'b1; //3
		14'b01110011001111: Borde = 1'b1; //4
		14'b01111011010000: Borde = 1'b1; //5
		14'b10000011010001: Borde = 1'b1; //6
		14'b10001011010010: Borde = 1'b1; //7
		
		14'b01010011101010: Borde = 1'b1; // 8
		14'b01011011101011: Borde = 1'b1; //9
		14'b01100011101100: Borde = 1'b1; //A
		14'b01101011101101: Borde = 1'b1; //B
		14'b01110011100101: Borde = 1'b1; // C
		14'b01111011100110: Borde = 1'b1; // D
		14'b10000011100111: Borde = 1'b1; // E
		14'b10001011101000: Borde = 1'b1; //F
		14'b10010011100100: Borde = 1'b1;// =
		
		14'b01010100011001: Borde = 1'b1; // punto
		14'b01011100001001: Borde = 1'b1; // raiz
		14'b01100100000010: Borde = 1'b1;//x
		14'b01101100000011: Borde = 1'b1;//division
		14'b01110100000000: Borde = 1'b1;//+
		14'b01111100000001: Borde = 1'b1;//-
		14'b10000100010011: Borde = 1'b1; // AC
		14'b10001100001110: Borde = 1'b1; // Borrar <-
		14'b10010100011000: Borde = 1'b1; // C borrar
		
	
		default: Borde = 1'b0;
	endcase
endmodule

//			1: Pos = 5'd20;		//0
//			2: Pos = 5'd21;		//1
//			4: Pos = 5'd22;		//2
//			8: Pos = 5'd23;		//3
//			16: Pos = 5'd15;		//4
//			32: Pos = 5'd16;		//5
//			64: Pos = 5'd17;		//6
//			128: Pos = 5'd18;		//7
//			256: Pos = 5'd10;		//8
//			512: Pos = 5'd11;		//9
//			1024: Pos = 5'd12;	//A
//			2048: Pos = 5'd13;	//B
//			4096: Pos = 5'd5;		//C
//			8192: Pos = 5'd6;		//D
//			16384: Pos = 5'd7;		//E
//			32768: Pos = 5'd8;		//F
//			65536: Pos = 5'd25;	// .  punto
//			131072: Pos = 5'd9;		//RAIZ
//			262144: Pos = 5'd2;		// X
//			524288: Pos = 5'd3;		// /
//			1048576: Pos = 5'd0;		// +
//			2097152: Pos = 5'd1;		// -
//			4194304: Pos = 5'd19;		//AC
//			8388608: Pos = 5'd14;		//BORRAR
//			16777216: Pos = 5'd24;		//CE delete
//			33554432: Pos = 5'd4;		// =
//			default: Pos = 5'd20;			//DEFAULT 0





//    3'b01000100000000: Borde = 1'b1;
//		3'b01001100000001: Borde = 1'b1;
//		3'b01010100000010: Borde = 1'b1;
//		3'b01011100000011: Borde = 1'b1;
//		3'b01100100000100: Borde = 1'b1;
//		
//		3'b01000100100101: Borde = 1'b1;
//		3'b01001100100110: Borde = 1'b1;
//		3'b01010100100111: Borde = 1'b1;
//		3'b01011100101000: Borde = 1'b1;
//		3'b01100100101001: Borde = 1'b1;
//		
//		3'b01000101001010: Borde = 1'b1;
//		3'b01001101001011: Borde = 1'b1;
//		3'b01010101001100: Borde = 1'b1;
//		3'b01011101001101: Borde = 1'b1;
//		3'b01100101001110: Borde = 1'b1;
//		
//		3'b01000101101111: Borde = 1'b1;
//		3'b01001101110000: Borde = 1'b1;
//		3'b01010101110001: Borde = 1'b1;
//		3'b01011101110010: Borde = 1'b1;
//		3'b01100101110011: Borde = 1'b1;
//		
//		3'b01000110010100: Borde = 1'b1;
//		3'b01001110010101: Borde = 1'b1;
//		3'b01010110010110: Borde = 1'b1;
//		3'b01011110010111: Borde = 1'b1;
//		3'b01100110011000: Borde = 1'b1;