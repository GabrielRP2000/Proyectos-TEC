`timescale 1ns / 1ps

module RomRegRotate16bits(SEL,WR);
	input [3:0] SEL;
	output reg [15:0] WR;

	always @(SEL)
		case (SEL)
			4'b0000: WR={4'b0000,4'b0000,4'b0000,4'b0001};
			4'b0001: WR={4'b0000,4'b0000,4'b0000,4'b0010};
			4'b0010: WR={4'b0000,4'b0000,4'b0000,4'b0100};
			4'b0011: WR={4'b0000,4'b0000,4'b0000,4'b1000};
			
			4'b0100: WR={4'b0000,4'b0000,4'b0001,4'b0000};
			4'b0101: WR={4'b0000,4'b0000,4'b0010,4'b0000};
			4'b0110: WR={4'b0000,4'b0000,4'b0100,4'b0000};
			4'b0111: WR={4'b0000,4'b0000,4'b1000,4'b0000};
			
			4'b1000: WR={4'b0000,4'b0001,4'b0000,4'b0000};
			4'b1001: WR={4'b0000,4'b0010,4'b0000,4'b0000};
			4'b1010: WR={4'b0000,4'b0100,4'b0000,4'b0000};
			4'b1011: WR={4'b0000,4'b1000,4'b0000,4'b0000};
			
			4'b1100: WR={4'b0001,4'b0000,4'b0000,4'b0000};
			4'b1101: WR={4'b0010,4'b0000,4'b0000,4'b0000};
			4'b1110: WR={4'b0100,4'b0000,4'b0000,4'b0000};
			4'b1111: WR={4'b1000,4'b0000,4'b0000,4'b0000};
	endcase
	
endmodule
